Current mirror sample
mp1 net01 net01 net11 vdd PMOS L=1.5u W=4u
mp2 net02 net01 net21 vdd PMOS L=1.5u W=4u

mp11 net11 vdd net12 vdd PMOS
mp12 net12 vdd net13 vdd PMOS
mp13 net13 vdd net14 vdd PMOS
mp14 net14 vdd vdd vdd PMOS
mp21 net21 vdd net22 vdd PMOS
mp22 net22 vdd net23 vdd PMOS
mp23 net23 vdd net24 vdd PMOS
mp24 net24 vdd vdd vdd PMOS

mp3 vout net02 vdd vdd PMOS L=1.5u W=4u
mn1 net11 gnd net04 gnd NMOS L=1.5u W=4u
mn2 net02 gnd net04 gnd NMOS L=1.5u W=4u
mn3 net05 net05 gnd gnd NMOS L=1.5u W=4u
mn4 net04 net05 gnd gnd NMOS L=1.5u W=4u
mn5 vout net05 gnd gnd NMOS L=1.5u W=4u

.MODEL PMOS pmos (VTO=-0.8V KP=5e-4 LAMBDA=0.01)

.MODEL NMOS nmos (VTO=-0.8V KP=5e-4 LAMBDA=0.01)

.AC dec 10 .01 10
.DC vs 0 5 0.05
.PROBE
.END
